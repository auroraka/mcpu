library verilog;
use verilog.vl_types.all;
entity rom_tf is
end rom_tf;
